// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Aug 16 14:45:23 2023"

module Zero(
	Zero
);


output wire	[31:0] Zero;

wire	[31:0] Zero_ALTERA_SYNTHESIZED;




































assign	Zero = Zero_ALTERA_SYNTHESIZED;
assign	Zero_ALTERA_SYNTHESIZED[0] = 0;
assign	Zero_ALTERA_SYNTHESIZED[1] = 0;
assign	Zero_ALTERA_SYNTHESIZED[2] = 0;
assign	Zero_ALTERA_SYNTHESIZED[3] = 0;
assign	Zero_ALTERA_SYNTHESIZED[4] = 0;
assign	Zero_ALTERA_SYNTHESIZED[5] = 0;
assign	Zero_ALTERA_SYNTHESIZED[6] = 0;
assign	Zero_ALTERA_SYNTHESIZED[7] = 0;
assign	Zero_ALTERA_SYNTHESIZED[8] = 0;
assign	Zero_ALTERA_SYNTHESIZED[9] = 0;
assign	Zero_ALTERA_SYNTHESIZED[10] = 0;
assign	Zero_ALTERA_SYNTHESIZED[11] = 0;
assign	Zero_ALTERA_SYNTHESIZED[12] = 0;
assign	Zero_ALTERA_SYNTHESIZED[13] = 0;
assign	Zero_ALTERA_SYNTHESIZED[14] = 0;
assign	Zero_ALTERA_SYNTHESIZED[15] = 0;
assign	Zero_ALTERA_SYNTHESIZED[16] = 0;
assign	Zero_ALTERA_SYNTHESIZED[31] = 0;
assign	Zero_ALTERA_SYNTHESIZED[30] = 0;
assign	Zero_ALTERA_SYNTHESIZED[29] = 0;
assign	Zero_ALTERA_SYNTHESIZED[28] = 0;
assign	Zero_ALTERA_SYNTHESIZED[27] = 0;
assign	Zero_ALTERA_SYNTHESIZED[26] = 0;
assign	Zero_ALTERA_SYNTHESIZED[25] = 0;
assign	Zero_ALTERA_SYNTHESIZED[24] = 0;
assign	Zero_ALTERA_SYNTHESIZED[23] = 0;
assign	Zero_ALTERA_SYNTHESIZED[22] = 0;
assign	Zero_ALTERA_SYNTHESIZED[21] = 0;
assign	Zero_ALTERA_SYNTHESIZED[20] = 0;
assign	Zero_ALTERA_SYNTHESIZED[19] = 0;
assign	Zero_ALTERA_SYNTHESIZED[18] = 0;
assign	Zero_ALTERA_SYNTHESIZED[17] = 0;

endmodule
